module alu_risc(

); 
endmodule


