module test(
	input a,
	input b,
	output c

),

endmodule